//-----------------------------------------------------------------------------
//
// Title       : test_Register
// Design      : DSD_Project
// Author      : shimu
// Company     : hp
//
//-----------------------------------------------------------------------------
//
// File        : C:/Users/HP/Downloads/DSD_Project/DSD_Project/DSD_Project/src/test_Register.v
// Generated   : Mon Jan 20 00:26:42 2025
// From        : Interface description file
// By          : ItfToHdl ver. 1.0
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------

`timescale 1ps / 1ps

//{{ Section below this comment is automatically maintained
//    and may be overwritten
//{module {test_Register}}

module test_Register ();

//}} End of automatically maintained section

// Enter your statements here //

endmodule
